-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 07 18:54:13 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MicroMouse IS
    PORT (
        reset : IN STD_LOGIC;
        clock : IN STD_LOGIC;
        Izquierda : IN STD_LOGIC;
        Derecha : IN STD_LOGIC;
        MI0 : OUT STD_LOGIC;
        MI1 : OUT STD_LOGIC;
        MD0 : OUT STD_LOGIC;
        MD1 : OUT STD_LOGIC
 );
END MicroMouse;

ARCHITECTURE BEHAVIOR OF MicroMouse IS
    TYPE type_fstate IS (stop,derecha90,izquierda90,giro180);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_MI0 : STD_LOGIC := '0';
    SIGNAL reg_MI1 : STD_LOGIC := '0';
    SIGNAL reg_MD0 : STD_LOGIC := '0';
    SIGNAL reg_MD1 : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
		  if reset = '0' then
				fstate <= stop;
        elsIF (RISING_EDGE(clock)) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Izquierda,Derecha,reg_MI0,reg_MI1,reg_MD0,reg_MD1)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= stop;
            reg_MI0 <= '0';
            reg_MI1 <= '0';
            reg_MD0 <= '0';
            reg_MD1 <= '0';
            MI0 <= '0';
            MI1 <= '0';
            MD0 <= '0';
            MD1 <= '0';
        ELSE
            reg_MI0 <= '0';
            reg_MI1 <= '0';
            reg_MD0 <= '0';
            reg_MD1 <= '0';
            MI0 <= '0';
            MI1 <= '0';
            MD0 <= '0';
            MD1 <= '0';
            CASE fstate IS
                WHEN stop =>
                    IF (((Izquierda = '0') AND (Derecha = '1'))) THEN
                        reg_fstate <= derecha90;
                    ELSIF (((Izquierda = '1') AND (Derecha = '0'))) THEN
                        reg_fstate <= izquierda90;
                    ELSIF (((Izquierda = '0') AND (Derecha = '0'))) THEN
                        reg_fstate <= stop;
                    ELSIF (((Izquierda = '1') AND (Derecha = '1'))) THEN
                        reg_fstate <= giro180;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= stop;
                    END IF;

                    reg_MI1 <= '0';

                    reg_MI0 <= '0';

                    reg_MD1 <= '0';

                    reg_MD0 <= '0';
                WHEN derecha90 =>
                    IF (((Izquierda = '0') AND (Derecha = '0'))) THEN
                        reg_fstate <= stop;
                    ELSIF (((Izquierda = '1') AND (Derecha = '1'))) THEN
                        reg_fstate <= giro180;
                    ELSIF (((Izquierda = '0') AND (Derecha = '1'))) THEN
                        reg_fstate <= derecha90;
                    ELSIF (((Izquierda = '1') AND (Derecha = '0'))) THEN
                        reg_fstate <= izquierda90;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= derecha90;
                    END IF;

						  reg_MI0 <= '1';
						  
                    reg_MI1 <= '0';

                    reg_MD0 <= '1';

                    reg_MD1 <= '0';
						  
                WHEN izquierda90 =>
                    IF (((Izquierda = '1') AND (Derecha = '1'))) THEN
                        reg_fstate <= giro180;
                    ELSIF (((Izquierda = '0') AND (Derecha = '0'))) THEN
                        reg_fstate <= stop;
                    ELSIF (((Izquierda = '1') AND (Derecha = '0'))) THEN
                        reg_fstate <= izquierda90;
                    ELSIF (((Izquierda = '0') AND (Derecha = '1'))) THEN
                        reg_fstate <= derecha90;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= izquierda90;
                    END IF;

                    reg_MI0 <= '0';

                    reg_MI1 <= '1';

                    reg_MD0 <= '0';

                    reg_MD1 <= '1';
                WHEN giro180 =>
                    IF (((Izquierda = '0') AND (Derecha = '0'))) THEN
                        reg_fstate <= stop;
                    ELSIF (((Izquierda = '0') AND (Derecha = '1'))) THEN
                        reg_fstate <= derecha90;
                    ELSIF (((Izquierda = '1') AND (Derecha = '0'))) THEN
                        reg_fstate <= izquierda90;
                    ELSIF (((Izquierda = '1') AND (Derecha = '1'))) THEN
                        reg_fstate <= giro180;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= giro180;
                    END IF;

						  reg_MI0 <= '1';
						  
                    reg_MI1 <= '0';

                    reg_MD0 <= '1';

                    reg_MD1 <= '0';
                WHEN OTHERS => 
                    reg_MI0 <= 'X';
                    reg_MI1 <= 'X';
                    reg_MD0 <= 'X';
                    reg_MD1 <= 'X';
                    report "Reach undefined state";
            END CASE;
            MI0 <= reg_MI0;
            MI1 <= reg_MI1;
            MD0 <= reg_MD0;
            MD1 <= reg_MD1;
        END IF;
    END PROCESS;
END BEHAVIOR;
